module InsMEM(
    input [31:0] addr,
    output reg [31:0] out
);
always@(addr)begin
    case(addr)
			32'd0:
				out <= 32'b1110_00_1_1101_0_0000_0000_000000010100;
			32'd8:
				out <= 32'b1110_00_1_1101_0_0000_0001_101000000001; 
			32'd8:
				out <= 32'b1110_00_1_1101_0_0000_0010_000100000011;
			32'd12:
				out <= 32'b1110_00_0_0100_1_0010_0011_000000000010;
			32'd16:
				out <= 32'b1110_00_0_0101_0_0000_0100_000000000000;
			32'd20:
				out <= 32'b1110_00_0_0010_0_0100_0101_000100000100;
			32'd24:
				out <= 32'b1110_00_0_0110_0_0000_0110_000010100000;
			32'd28:
				out <= 32'b1110_00_0_1100_0_0101_0111_000101000010; 
			32'd32:
				out <= 32'b1110_00_0_0000_0_0111_1000_000000000011;
			32'd36:
				out <= 32'b1110_00_0_1111_0_0000_1001_000000000110;
			32'd40:
				out <= 32'b1110_00_0_0001_0_0100_1010_000000000101;
			32'd44:
				out <= 32'b1110_00_0_1010_1_1000_0000_000000000110;
			32'd48:
				out <= 32'b0001_00_0_0100_0_0001_0001_000000000001; 
			32'd52:
				out <= 32'b1110_00_0_1000_1_1001_0000_000000001000; 
			32'd56:
				out <= 32'b0000_00_0_0100_0_0010_0010_000000000010;
			32'd60:
				out <= 32'b1110_00_1_1101_0_0000_0000_101100000001; 
			32'd64:
				out <= 32'b1110_01_0_0100_0_0000_0001_000000000000;  
			32'd68:
				out <= 32'b1110_01_0_0100_1_0000_1011_000000000000; 
		endcase
	end
endmodule