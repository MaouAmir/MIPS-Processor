`timescale 1ns/1ns

module IF_TB();





endmodule
